LIBRARY IEEE;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_4X1_NBITS IS
   GENERIC(
      N  : INTEGER := 4   -- Length of each signal input (X bits)
   );
   PORT(
      i_BUS_A   :   IN    STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_BUS_B   :   IN    STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_BUS_C   :   IN    STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_BUS_D   :   IN    STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_SEL     :   IN    STD_LOGIC_VECTOR( 1  DOWNTO 0);
      o_BUS     :   OUT   STD_LOGIC_VECTOR(N-1 DOWNTO 0)
   );
END MUX_4X1_NBITS;

ARCHITECTURE BEHAVIORAL OF MUX_4X1_NBITS IS
BEGIN
   WITH i_SEL SELECT
      o_BUS <= i_BUS_A WHEN "00",
      i_BUS_B WHEN "01",
      i_BUS_C WHEN "10",
      i_BUS_D WHEN "11",
   (OTHERS =>'Z') WHEN OTHERS;
END BEHAVIORAL;
