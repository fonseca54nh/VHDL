LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY HALF_SUBTRACTOR IS
PORT(
   i_A        :   IN    STD_LOGIC;
   i_B        :   IN    STD_LOGIC;
   o_Diff     :   OUT   STD_LOGIC;
   o_Borrow   :   OUT   STD_LOGIC
);
END HALF_SUBTRACTOR;

ARCHITECTURE STRUCTURAL OF HALF_SUBTRACTOR IS
BEGIN
   o_Diff   <= i_A XOR i_B;
   o_Borrow <= (NOT i_A) AND i_B;
END STRUCTURAL;
