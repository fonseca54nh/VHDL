LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY AND_GENERATE IS
   GENERIC(
      N      :   INTEGER := 16
   );
   PORT(
      i_A    :   IN   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_B    :   IN   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_C    :   IN   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_D    :   IN   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      i_E    :   IN   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
      o_C    :   OUT  STD_LOGIC_VECTOR(N-1 DOWNTO 0)
   );
END AND_GENERATE;

ARCHITECTURE BEHAVIORAL OF AND_GENERATE IS
   SIGNAL w_F   :   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
   SIGNAL w_G   :   STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN
   U01 : FOR i IN (N-1) DOWNTO 0 GENERATE
      w_F(i) <= i_A(i) AND i_B(i) AND i_C(i);
      w_G(i) <= i_C(i) AND i_D(i) AND i_E(i);
      o_C(i) <= w_F(i) OR  w_G(i);
   END GENERATE U01;	
END BEHAVIORAL;
