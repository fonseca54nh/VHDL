LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY FlipFlopAsync IS
	PORT (
		i_RST   :  IN   STD_LOGIC;
		i_CLK   :  IN   STD_LOGIC;
		i_DATA  :  IN   STD_LOGIC;
		o_DATA  :  out  STD_LOGIC
	);
END FlipFlopAsync;

ARCHITECTURE BEHAVIORAL OF FlipFlopAsync IS

BEGIN

	PROCESS(i_CLK, i_RST)
	BEGIN
		IF (i_RST = '1') THEN
			o_DATA <= '0';
		ELSE 	
			IF RISING_EDGE(i_CLK) THEN 
			   o_DATA <= i_DATA;
			END IF;
		END IF;
	END PROCESS;

END BEHAVIORAL;
